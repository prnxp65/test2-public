# Copyright (c) NXP Semiconductors
# NXP Confidential Proprietary
# Compiler: s10hv_1prf
# Revision: s10hv_1prf_1.11.01 
# Date: Sun Apr 03 20:50:56 MST 2022

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO s10hv_1prf_w1024x16b1c08_ulm
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN s10hv_1prf_w1024x16b1c08_ulm 0 0 ;
  SIZE 302.4 BY 342.72 ;
  SYMMETRY X Y R90 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.77675 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.88 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER m3 ;
      ANTENNAMAXAREACAR 22.157083 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 81.227778 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 108.21 0 108.51 0.68 ;
      LAYER m2 ;
        RECT 108.21 0 108.51 0.68 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.75025 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.7 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER m3 ;
      ANTENNAMAXAREACAR 17.073472 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 64.027778 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 110.73 0 111.03 0.68 ;
      LAYER m2 ;
        RECT 110.73 0 111.03 0.68 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.74165 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.396 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER m3 ;
      ANTENNAMAXAREACAR 17.034583 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 63.133333 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 113.25 0 113.55 0.68 ;
      LAYER m2 ;
        RECT 113.25 0 113.55 0.68 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8529 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.408 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER m3 ;
      ANTENNAMAXAREACAR 29.641389 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 109.719444 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 130.89 0 131.19 0.68 ;
      LAYER m2 ;
        RECT 130.89 0 131.19 0.68 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.729 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.936 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER m3 ;
      ANTENNAMAXAREACAR 29.626389 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 109.066667 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 140.97 0 141.27 0.68 ;
      LAYER m2 ;
        RECT 140.97 0 141.27 0.68 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.8655 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.456 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER m3 ;
      ANTENNAMAXAREACAR 29.561111 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 109.611111 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 166.17 0 166.47 0.68 ;
      LAYER m2 ;
        RECT 166.17 0 166.47 0.68 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.1574 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.568 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER m3 ;
      ANTENNAMAXAREACAR 31.955972 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 118.325 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 118.29 0 118.59 0.68 ;
      LAYER m2 ;
        RECT 118.29 0 118.59 0.68 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.86195 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER m3 ;
      ANTENNAMAXAREACAR 31.265972 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 112.902778 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 120.81 0 121.11 0.68 ;
      LAYER m2 ;
        RECT 120.81 0 121.11 0.68 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.79725 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.196 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER m3 ;
      ANTENNAMAXAREACAR 28.295139 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 106.747222 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 128.37 0 128.67 0.68 ;
      LAYER m2 ;
        RECT 128.37 0 128.67 0.68 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.88545 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 37.532 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.36 LAYER m3 ;
      ANTENNAMAXAREACAR 28.611528 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 108.188889 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 168.69 0 168.99 0.68 ;
      LAYER m2 ;
        RECT 168.69 0 168.99 0.68 ;
    END
  END a[9]
  PIN cen_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2698 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.52 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.45 LAYER m3 ;
      ANTENNAMAXAREACAR 16.014667 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 52.44 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 135.93 0 136.23 0.68 ;
      LAYER m2 ;
        RECT 135.93 0 136.23 0.68 ;
    END
  END cen_b
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5512 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.592 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 2.628 LAYER m3 ;
      ANTENNAMAXAREACAR 7.197807 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 21.736894 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 146.01 0 146.31 0.68 ;
      LAYER m2 ;
        RECT 146.01 0 146.31 0.68 ;
    END
  END clk
  PIN d[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 7.41 0 7.71 0.68 ;
      LAYER m2 ;
        RECT 7.41 0 7.71 0.68 ;
    END
  END d[0]
  PIN d[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 224.13 0 224.43 0.68 ;
      LAYER m2 ;
        RECT 224.13 0 224.43 0.68 ;
    END
  END d[10]
  PIN d[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.22545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.441 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.88642 LAYER m3 ;
      ANTENNAMAXAREACAR 5.25679 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 17.037037 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.222222 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 236.73 0 237.03 0.68 ;
      LAYER m2 ;
        RECT 236.73 0 237.03 0.68 ;
    END
  END d[11]
  PIN d[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 249.33 0 249.63 0.68 ;
      LAYER m2 ;
        RECT 249.33 0 249.63 0.68 ;
    END
  END d[12]
  PIN d[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 261.93 0 262.23 0.68 ;
      LAYER m2 ;
        RECT 261.93 0 262.23 0.68 ;
    END
  END d[13]
  PIN d[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 274.53 0 274.83 0.68 ;
      LAYER m2 ;
        RECT 274.53 0 274.83 0.68 ;
    END
  END d[14]
  PIN d[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 287.13 0 287.43 0.68 ;
      LAYER m2 ;
        RECT 287.13 0 287.43 0.68 ;
    END
  END d[15]
  PIN d[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 20.01 0 20.31 0.68 ;
      LAYER m2 ;
        RECT 20.01 0 20.31 0.68 ;
    END
  END d[1]
  PIN d[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 32.61 0 32.91 0.68 ;
      LAYER m2 ;
        RECT 32.61 0 32.91 0.68 ;
    END
  END d[2]
  PIN d[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 45.21 0 45.51 0.68 ;
      LAYER m2 ;
        RECT 45.21 0 45.51 0.68 ;
    END
  END d[3]
  PIN d[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 57.81 0 58.11 0.68 ;
      LAYER m2 ;
        RECT 57.81 0 58.11 0.68 ;
    END
  END d[4]
  PIN d[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 70.41 0 70.71 0.68 ;
      LAYER m2 ;
        RECT 70.41 0 70.71 0.68 ;
    END
  END d[5]
  PIN d[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 83.01 0 83.31 0.68 ;
      LAYER m2 ;
        RECT 83.01 0 83.31 0.68 ;
    END
  END d[6]
  PIN d[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 95.61 0 95.91 0.68 ;
      LAYER m2 ;
        RECT 95.61 0 95.91 0.68 ;
    END
  END d[7]
  PIN d[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 198.93 0 199.23 0.68 ;
      LAYER m2 ;
        RECT 198.93 0 199.23 0.68 ;
    END
  END d[8]
  PIN d[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.21545 LAYER m2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.411 LAYER m2 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324 LAYER m3 ;
      ANTENNAGATEAREA 0.324 LAYER m2 ;
      ANTENNAMAXAREACAR 5.855556 LAYER m3 ;
      ANTENNAMAXAREACAR 5.225926 LAYER m2 ;
      ANTENNAMAXSIDEAREACAR 16.944444 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 15.12963 LAYER m2 ;
      ANTENNAMAXCUTCAR 0.4 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 209.01 0 209.31 0.68 ;
      LAYER m2 ;
        RECT 209.01 0 209.31 0.68 ;
    END
  END d[9]
  PIN ipt_nowrite
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.96975 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.996 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.81 LAYER m3 ;
      ANTENNAMAXAREACAR 5.628889 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 20.969136 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 125.85 0 126.15 0.68 ;
      LAYER m2 ;
        RECT 125.85 0 126.15 0.68 ;
    END
  END ipt_nowrite
  PIN ipt_st_dis
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2051 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.896 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.45 LAYER m3 ;
      ANTENNAMAXAREACAR 11.688667 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 42.951111 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 133.41 0 133.71 0.68 ;
      LAYER m2 ;
        RECT 133.41 0 133.71 0.68 ;
    END
  END ipt_st_dis
  PIN q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 9.93 0 10.23 0.685 ;
      LAYER m2 ;
        RECT 9.93 0 10.23 0.685 ;
    END
  END q[0]
  PIN q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 226.65 0 226.95 0.685 ;
      LAYER m2 ;
        RECT 226.65 0 226.95 0.685 ;
    END
  END q[10]
  PIN q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 239.25 0 239.55 0.685 ;
      LAYER m2 ;
        RECT 239.25 0 239.55 0.685 ;
    END
  END q[11]
  PIN q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 251.85 0 252.15 0.685 ;
      LAYER m2 ;
        RECT 251.85 0 252.15 0.685 ;
    END
  END q[12]
  PIN q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 264.45 0 264.75 0.685 ;
      LAYER m2 ;
        RECT 264.45 0 264.75 0.685 ;
    END
  END q[13]
  PIN q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 277.05 0 277.35 0.685 ;
      LAYER m2 ;
        RECT 277.05 0 277.35 0.685 ;
    END
  END q[14]
  PIN q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 289.65 0 289.95 0.685 ;
      LAYER m2 ;
        RECT 289.65 0 289.95 0.685 ;
    END
  END q[15]
  PIN q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 22.53 0 22.83 0.685 ;
      LAYER m2 ;
        RECT 22.53 0 22.83 0.685 ;
    END
  END q[1]
  PIN q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 35.13 0 35.43 0.685 ;
      LAYER m2 ;
        RECT 35.13 0 35.43 0.685 ;
    END
  END q[2]
  PIN q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 47.73 0 48.03 0.685 ;
      LAYER m2 ;
        RECT 47.73 0 48.03 0.685 ;
    END
  END q[3]
  PIN q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 60.33 0 60.63 0.685 ;
      LAYER m2 ;
        RECT 60.33 0 60.63 0.685 ;
    END
  END q[4]
  PIN q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 72.93 0 73.23 0.685 ;
      LAYER m2 ;
        RECT 72.93 0 73.23 0.685 ;
    END
  END q[5]
  PIN q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 85.53 0 85.83 0.685 ;
      LAYER m2 ;
        RECT 85.53 0 85.83 0.685 ;
    END
  END q[6]
  PIN q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 98.13 0 98.43 0.685 ;
      LAYER m2 ;
        RECT 98.13 0 98.43 0.685 ;
    END
  END q[7]
  PIN q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 201.45 0 201.75 0.685 ;
      LAYER m2 ;
        RECT 201.45 0 201.75 0.685 ;
    END
  END q[8]
  PIN q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.73945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.304 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    PORT
      LAYER m3 ;
        RECT 214.05 0 214.35 0.685 ;
      LAYER m2 ;
        RECT 214.05 0 214.35 0.685 ;
    END
  END q[9]
  PIN valen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9238 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.44 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.375 LAYER m3 ;
      ANTENNAMAXAREACAR 17.3992 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 65.304 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 173.73 0 174.03 0.68 ;
      LAYER m2 ;
        RECT 173.73 0 174.03 0.68 ;
    END
  END valen
  PIN valrd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.09945 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.236 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER m3 ;
      ANTENNAMAXAREACAR 26.030426 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 95.375969 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 176.25 0 176.55 0.68 ;
      LAYER m2 ;
        RECT 176.25 0 176.55 0.68 ;
    END
  END valrd[0]
  PIN valrd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.8578 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.312 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER m3 ;
      ANTENNAMAXAREACAR 24.529457 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 91.189922 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 178.77 0 179.07 0.68 ;
      LAYER m2 ;
        RECT 178.77 0 179.07 0.68 ;
    END
  END valrd[1]
  PIN valrd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.90085 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.476 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER m3 ;
      ANTENNAMAXAREACAR 24.034302 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 91.116279 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 186.33 0 186.63 0.68 ;
      LAYER m2 ;
        RECT 186.33 0 186.63 0.68 ;
    END
  END valrd[2]
  PIN valwr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1971 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.608 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER m3 ;
      ANTENNAMAXAREACAR 25.182558 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 95.503876 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 188.85 0 189.15 0.68 ;
      LAYER m2 ;
        RECT 188.85 0 189.15 0.68 ;
    END
  END valwr[0]
  PIN valwr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.59635 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.316 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER m3 ;
      ANTENNAMAXAREACAR 22.85407 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 86.620155 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 191.37 0 191.67 0.68 ;
      LAYER m2 ;
        RECT 191.37 0 191.67 0.68 ;
    END
  END valwr[1]
  PIN valwr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6562 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.544 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.258 LAYER m3 ;
      ANTENNAMAXAREACAR 23.227132 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 87.655039 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 193.89 0 194.19 0.68 ;
      LAYER m2 ;
        RECT 193.89 0 194.19 0.68 ;
    END
  END valwr[2]
  PIN wen
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3416 LAYER m3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.416 LAYER m3 ;
    ANTENNAPARTIALCUTAREA 0.0648 LAYER via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.54 LAYER m3 ;
      ANTENNAMAXAREACAR 9.437963 LAYER m3 ;
      ANTENNAMAXSIDEAREACAR 34.95 LAYER m3 ;
    PORT
      LAYER m3 ;
        RECT 123.33 0 123.63 0.68 ;
      LAYER m2 ;
        RECT 123.33 0 123.63 0.68 ;
    END
  END wen
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER ulm ;
        RECT 0 323.83 302.4 328.84 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 307.99 302.4 313 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 292.15 302.4 297.16 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 276.31 302.4 281.32 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 260.47 302.4 265.48 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 244.63 302.4 249.64 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 228.79 302.4 233.8 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 212.95 302.4 217.96 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 197.11 302.4 202.12 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 181.27 302.4 186.28 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 165.43 302.4 170.44 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 149.59 302.4 154.6 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 133.75 302.4 138.76 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 117.91 302.4 122.92 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 102.07 302.4 107.08 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 86.23 302.4 91.24 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 71.04 302.4 76.05 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 39.58 302.4 44.59 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 19.06 302.4 24.07 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER ulm ;
        RECT 0 331.75 302.4 336.76 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 315.91 302.4 320.92 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 300.07 302.4 305.08 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 284.23 302.4 289.24 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 268.39 302.4 273.4 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 252.55 302.4 257.56 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 236.71 302.4 241.72 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 220.87 302.4 225.88 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 205.03 302.4 210.04 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 189.19 302.4 194.2 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 173.35 302.4 178.36 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 157.51 302.4 162.52 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 141.67 302.4 146.68 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 125.83 302.4 130.84 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 109.99 302.4 115 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 94.15 302.4 99.16 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 78.31 302.4 83.32 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 32.57 302.4 37.58 ;
    END
    PORT
      LAYER ulm ;
        RECT 0 12.05 302.4 17.06 ;
    END
  END vss
  OBS
    LAYER m3 ;
      RECT 191.03 27.665 191.33 78.355 ;
      RECT 191.03 27.665 192.005 27.965 ;
      RECT 191.705 1.275 192.005 27.965 ;
      RECT 182.415 0.48 182.625 5.115 ;
      RECT 182.415 0.48 184.11 0.69 ;
      RECT 183.81 0 184.11 0.69 ;
      RECT 181.29 0 181.5 5.115 ;
      RECT 181.29 0 181.59 0.68 ;
      RECT 115.815 0 116.025 5.115 ;
      RECT 115.77 0 116.07 0.68 ;
      RECT 297.86 2.56 298.16 78.055 ;
      RECT 297.2 2.56 297.5 78.055 ;
      RECT 288.675 4.015 288.885 8.25 ;
      RECT 276.915 4.015 277.125 8.25 ;
      RECT 272.96 2.56 273.26 78.055 ;
      RECT 272.3 2.56 272.66 78.055 ;
      RECT 271.7 2.56 272 78.055 ;
      RECT 263.175 4.015 263.385 8.25 ;
      RECT 251.415 4.015 251.625 8.25 ;
      RECT 247.46 2.56 247.76 78.055 ;
      RECT 246.8 2.56 247.16 78.055 ;
      RECT 246.2 2.56 246.5 78.055 ;
      RECT 237.675 4.015 237.885 8.25 ;
      RECT 225.915 4.015 226.125 8.25 ;
      RECT 221.96 2.56 222.26 78.055 ;
      RECT 221.3 2.56 221.66 78.055 ;
      RECT 220.7 2.56 221 78.055 ;
      RECT 217.445 3.66 217.655 13.32 ;
      RECT 212.175 4.015 212.385 8.25 ;
      RECT 205.685 3.66 205.895 13.32 ;
      RECT 200.415 4.015 200.625 8.25 ;
      RECT 196.46 2.56 196.76 78.055 ;
      RECT 195.8 2.56 196.16 78.055 ;
      RECT 195.2 2.56 195.5 78.055 ;
      RECT 194.44 4.01 194.65 5.145 ;
      RECT 191.195 4.01 191.405 5.14 ;
      RECT 190.37 1.275 190.67 78.355 ;
      RECT 186.38 2.52 187.04 78.055 ;
      RECT 185.855 4.01 186.065 5.785 ;
      RECT 185.01 4.01 185.22 5.16 ;
      RECT 183.425 1.275 184.085 78.055 ;
      RECT 180.28 4.01 180.49 5.325 ;
      RECT 179.35 1.275 180.01 45.075 ;
      RECT 178.87 4.01 179.08 5.505 ;
      RECT 177.305 2.525 177.965 78.055 ;
      RECT 175.21 1.275 175.87 44.76 ;
      RECT 174.495 4.01 174.705 5.115 ;
      RECT 171.2 1.275 171.86 47.515 ;
      RECT 169.84 4.01 170.05 5.115 ;
      RECT 167.96 1.275 168.62 47.515 ;
      RECT 167.3 4.01 167.51 5.115 ;
      RECT 164.735 1.275 165.395 78.055 ;
      RECT 161.365 1.275 162.025 78.055 ;
      RECT 158.225 1.275 158.885 78.055 ;
      RECT 156.62 1.275 157.28 47.515 ;
      RECT 154.79 1.275 155.45 45.075 ;
      RECT 145.335 4.01 145.545 5.115 ;
      RECT 142.02 1.275 142.68 45.075 ;
      RECT 141.375 4.01 141.585 5.115 ;
      RECT 140.19 1.275 140.85 47.515 ;
      RECT 138.585 1.275 139.245 78.055 ;
      RECT 135.445 1.275 136.105 78.055 ;
      RECT 134.535 4.01 134.745 5.115 ;
      RECT 132.075 2.52 132.735 78.055 ;
      RECT 131.295 4.01 131.505 5.925 ;
      RECT 130.215 4.01 130.425 5.115 ;
      RECT 128.85 1.275 129.51 47.515 ;
      RECT 127.695 4.01 127.905 5.115 ;
      RECT 125.61 1.275 126.27 47.515 ;
      RECT 124.815 4.01 125.025 5.115 ;
      RECT 121.6 2.555 122.26 45.075 ;
      RECT 120.855 4.01 121.065 5.875 ;
      RECT 119.505 2.54 120.165 78.055 ;
      RECT 118.695 4.01 118.905 6.075 ;
      RECT 117.46 1.275 118.12 45.075 ;
      RECT 116.895 4.01 117.105 5.115 ;
      RECT 114.735 4.01 114.945 5.115 ;
      RECT 113.385 1.275 114.045 78.055 ;
      RECT 112.575 4.01 112.785 5.115 ;
      RECT 111.495 4.01 111.705 6.09 ;
      RECT 110.43 2.52 111.09 78.055 ;
      RECT 106.8 2.56 107.1 78.055 ;
      RECT 106.14 2.56 106.44 78.055 ;
      RECT 97.615 4.015 97.825 8.25 ;
      RECT 85.855 4.015 86.065 8.25 ;
      RECT 81.9 2.56 82.2 78.055 ;
      RECT 81.24 2.56 81.6 78.055 ;
      RECT 80.64 2.56 80.94 78.055 ;
      RECT 72.115 4.015 72.325 8.25 ;
      RECT 60.355 4.015 60.565 8.25 ;
      RECT 56.4 2.56 56.7 78.055 ;
      RECT 55.74 2.56 56.1 78.055 ;
      RECT 55.14 2.56 55.44 78.055 ;
      RECT 46.615 4.015 46.825 8.25 ;
      RECT 34.855 4.015 35.065 8.25 ;
      RECT 30.9 2.56 31.2 78.055 ;
      RECT 30.24 2.56 30.6 78.055 ;
      RECT 29.64 2.56 29.94 78.055 ;
      RECT 21.115 4.015 21.325 8.25 ;
      RECT 9.355 4.015 9.565 8.25 ;
      RECT 5.4 2.56 5.7 78.055 ;
      RECT 4.74 2.56 5.04 78.055 ;
    LAYER m3 SPACING 0.21 ;
      RECT 0 0.895 302.4 342.72 ;
      RECT 290.16 0 302.4 342.72 ;
      RECT 277.56 0.89 289.44 342.72 ;
      RECT 287.64 0 289.44 342.72 ;
      RECT 264.96 0.89 276.84 342.72 ;
      RECT 275.04 0 276.84 342.72 ;
      RECT 252.36 0.89 264.24 342.72 ;
      RECT 262.44 0 264.24 342.72 ;
      RECT 239.76 0.89 251.64 342.72 ;
      RECT 249.84 0 251.64 342.72 ;
      RECT 227.16 0.89 239.04 342.72 ;
      RECT 237.24 0 239.04 342.72 ;
      RECT 214.56 0.89 226.44 342.72 ;
      RECT 224.64 0 226.44 342.72 ;
      RECT 201.96 0.89 213.84 342.72 ;
      RECT 209.52 0 213.84 342.72 ;
      RECT 98.64 0.89 201.24 342.72 ;
      RECT 199.44 0 201.24 342.72 ;
      RECT 86.04 0.89 97.92 342.72 ;
      RECT 96.12 0 97.92 342.72 ;
      RECT 73.44 0.89 85.32 342.72 ;
      RECT 83.52 0 85.32 342.72 ;
      RECT 60.84 0.89 72.72 342.72 ;
      RECT 70.92 0 72.72 342.72 ;
      RECT 48.24 0.89 60.12 342.72 ;
      RECT 58.32 0 60.12 342.72 ;
      RECT 35.64 0.89 47.52 342.72 ;
      RECT 45.72 0 47.52 342.72 ;
      RECT 23.04 0.89 34.92 342.72 ;
      RECT 33.12 0 34.92 342.72 ;
      RECT 10.44 0.89 22.32 342.72 ;
      RECT 20.52 0 22.32 342.72 ;
      RECT 0 0.89 9.72 342.72 ;
      RECT 7.92 0 9.72 342.72 ;
      RECT 277.56 0 286.92 342.72 ;
      RECT 264.96 0 274.32 342.72 ;
      RECT 252.36 0 261.72 342.72 ;
      RECT 239.76 0 249.12 342.72 ;
      RECT 227.16 0 236.52 342.72 ;
      RECT 214.56 0 223.92 342.72 ;
      RECT 201.96 0 208.8 342.72 ;
      RECT 194.4 0 198.72 342.72 ;
      RECT 191.88 0 193.68 342.72 ;
      RECT 189.36 0 191.16 342.72 ;
      RECT 186.84 0 188.64 342.72 ;
      RECT 179.28 0 186.12 342.72 ;
      RECT 176.76 0 178.56 342.72 ;
      RECT 174.24 0 176.04 342.72 ;
      RECT 169.2 0 173.52 342.72 ;
      RECT 166.68 0 168.48 342.72 ;
      RECT 146.52 0 165.96 342.72 ;
      RECT 141.48 0 145.8 342.72 ;
      RECT 136.44 0 140.76 342.72 ;
      RECT 133.92 0 135.72 342.72 ;
      RECT 131.4 0 133.2 342.72 ;
      RECT 128.88 0 130.68 342.72 ;
      RECT 126.36 0 128.16 342.72 ;
      RECT 123.84 0 125.64 342.72 ;
      RECT 121.32 0 123.12 342.72 ;
      RECT 118.8 0 120.6 342.72 ;
      RECT 113.76 0 118.08 342.72 ;
      RECT 111.24 0 113.04 342.72 ;
      RECT 108.72 0 110.52 342.72 ;
      RECT 98.64 0 108 342.72 ;
      RECT 86.04 0 95.4 342.72 ;
      RECT 73.44 0 82.8 342.72 ;
      RECT 60.84 0 70.2 342.72 ;
      RECT 48.24 0 57.6 342.72 ;
      RECT 35.64 0 45 342.72 ;
      RECT 23.04 0 32.4 342.72 ;
      RECT 10.44 0 19.8 342.72 ;
      RECT 0 0 7.2 342.72 ;
    LAYER m2 ;
      RECT 211.185 0.86 211.395 3.435 ;
      RECT 210.915 0.86 211.48 1.07 ;
      RECT 84.865 2.285 85.075 3.435 ;
      RECT 84.915 0.86 85.075 3.435 ;
      RECT 84.915 0.86 85.16 1.07 ;
      RECT 296.99 4.31 301.845 4.97 ;
      RECT 296.99 6.585 301.845 7.245 ;
      RECT 296.99 8.515 301.845 9.175 ;
      RECT 296.99 11.42 301.845 12.08 ;
      RECT 296.99 14.485 301.845 15.025 ;
      RECT 296.99 17.725 301.845 18.265 ;
      RECT 296.99 23.555 301.845 24.095 ;
      RECT 296.99 25.7 301.845 26.24 ;
      RECT 296.99 27.86 301.845 28.4 ;
      RECT 296.99 30.755 301.845 31.295 ;
      RECT 296.99 32.98 301.845 33.52 ;
      RECT 296.99 34.475 301.845 35.015 ;
      RECT 296.99 36.895 301.845 37.435 ;
      RECT 296.99 37.675 301.845 38.335 ;
      RECT 296.99 42.835 301.845 43.495 ;
      RECT 297.2 52.49 301.845 53.03 ;
      RECT 296.99 54.05 301.845 54.53 ;
      RECT 296.99 55.28 301.845 55.76 ;
      RECT 297.2 56.78 301.845 57.32 ;
      RECT 296.99 66.37 301.845 66.91 ;
      RECT 296.99 69.65 301.845 70.98 ;
      RECT 296.99 72.95 301.845 74.28 ;
      RECT 296.99 74.995 301.845 75.655 ;
      RECT 296.99 76.8 301.845 77.46 ;
      RECT 287.685 2.285 287.895 3.435 ;
      RECT 285.38 0.86 285.525 1.07 ;
      RECT 275.925 2.285 276.135 3.435 ;
      RECT 262.185 2.285 262.395 3.435 ;
      RECT 259.88 0.86 260.325 1.07 ;
      RECT 250.425 2.285 250.635 3.435 ;
      RECT 236.685 2.285 236.895 3.435 ;
      RECT 234.38 0.86 235.125 1.07 ;
      RECT 224.925 2.285 225.135 3.435 ;
      RECT 199.425 2.285 199.635 3.435 ;
      RECT 197.12 0.86 197.325 1.07 ;
      RECT 183.81 0 184.11 0.68 ;
      RECT 181.29 0 181.59 0.68 ;
      RECT 115.77 0 116.07 0.68 ;
      RECT 96.625 2.285 96.835 3.435 ;
      RECT 71.125 2.285 71.335 3.435 ;
      RECT 59.365 2.285 59.575 3.435 ;
      RECT 45.625 2.285 45.835 3.435 ;
      RECT 43.32 0.86 43.605 1.07 ;
      RECT 33.865 2.285 34.075 3.435 ;
      RECT 20.125 2.285 20.335 3.435 ;
      RECT 17.82 0.86 18.405 1.07 ;
      RECT 8.365 2.285 8.575 3.435 ;
      RECT 1.055 4.31 5.91 4.97 ;
      RECT 1.055 6.585 5.91 7.245 ;
      RECT 1.055 8.515 5.91 9.175 ;
      RECT 1.055 11.42 5.91 12.08 ;
      RECT 1.055 14.485 5.91 15.025 ;
      RECT 1.055 17.725 5.91 18.265 ;
      RECT 1.055 23.555 5.91 24.095 ;
      RECT 1.055 25.7 5.91 26.24 ;
      RECT 1.055 27.86 5.91 28.4 ;
      RECT 1.055 30.755 5.91 31.295 ;
      RECT 1.055 32.98 5.91 33.52 ;
      RECT 1.055 34.475 5.91 35.015 ;
      RECT 1.055 36.895 5.91 37.435 ;
      RECT 1.055 37.675 5.91 38.335 ;
      RECT 1.055 42.835 5.91 43.495 ;
      RECT 1.055 54.05 5.91 54.53 ;
      RECT 1.055 55.28 5.91 55.76 ;
      RECT 1.055 66.37 5.91 66.91 ;
      RECT 1.055 69.655 5.91 70.975 ;
      RECT 1.055 72.955 5.91 74.275 ;
      RECT 1.055 74.995 5.91 75.655 ;
      RECT 1.055 76.8 5.91 77.46 ;
      RECT 1.055 52.52 5.7 53 ;
      RECT 1.055 56.81 5.7 57.29 ;
    LAYER m2 SPACING 0.18 ;
      RECT 0 0.865 302.4 342.72 ;
      RECT 290.13 0 302.4 342.72 ;
      RECT 277.53 0.86 289.47 342.72 ;
      RECT 287.61 0 289.47 342.72 ;
      RECT 264.93 0.86 276.87 342.72 ;
      RECT 275.01 0 276.87 342.72 ;
      RECT 252.33 0.86 264.27 342.72 ;
      RECT 262.41 0 264.27 342.72 ;
      RECT 239.73 0.86 251.67 342.72 ;
      RECT 249.81 0 251.67 342.72 ;
      RECT 227.13 0.86 239.07 342.72 ;
      RECT 237.21 0 239.07 342.72 ;
      RECT 214.53 0.86 226.47 342.72 ;
      RECT 224.61 0 226.47 342.72 ;
      RECT 201.93 0.86 213.87 342.72 ;
      RECT 209.49 0 213.87 342.72 ;
      RECT 98.61 0.86 201.27 342.72 ;
      RECT 199.41 0 201.27 342.72 ;
      RECT 86.01 0.86 97.95 342.72 ;
      RECT 96.09 0 97.95 342.72 ;
      RECT 73.41 0.86 85.35 342.72 ;
      RECT 83.49 0 85.35 342.72 ;
      RECT 60.81 0.86 72.75 342.72 ;
      RECT 70.89 0 72.75 342.72 ;
      RECT 48.21 0.86 60.15 342.72 ;
      RECT 58.29 0 60.15 342.72 ;
      RECT 35.61 0.86 47.55 342.72 ;
      RECT 45.69 0 47.55 342.72 ;
      RECT 23.01 0.86 34.95 342.72 ;
      RECT 33.09 0 34.95 342.72 ;
      RECT 10.41 0.86 22.35 342.72 ;
      RECT 20.49 0 22.35 342.72 ;
      RECT 0 0.86 9.75 342.72 ;
      RECT 7.89 0 9.75 342.72 ;
      RECT 277.53 0 286.95 342.72 ;
      RECT 264.93 0 274.35 342.72 ;
      RECT 252.33 0 261.75 342.72 ;
      RECT 239.73 0 249.15 342.72 ;
      RECT 227.13 0 236.55 342.72 ;
      RECT 214.53 0 223.95 342.72 ;
      RECT 201.93 0 208.83 342.72 ;
      RECT 194.37 0 198.75 342.72 ;
      RECT 191.85 0 193.71 342.72 ;
      RECT 189.33 0 191.19 342.72 ;
      RECT 186.81 0 188.67 342.72 ;
      RECT 179.25 0 186.15 342.72 ;
      RECT 176.73 0 178.59 342.72 ;
      RECT 174.21 0 176.07 342.72 ;
      RECT 169.17 0 173.55 342.72 ;
      RECT 166.65 0 168.51 342.72 ;
      RECT 146.49 0 165.99 342.72 ;
      RECT 141.45 0 145.83 342.72 ;
      RECT 136.41 0 140.79 342.72 ;
      RECT 133.89 0 135.75 342.72 ;
      RECT 131.37 0 133.23 342.72 ;
      RECT 128.85 0 130.71 342.72 ;
      RECT 126.33 0 128.19 342.72 ;
      RECT 123.81 0 125.67 342.72 ;
      RECT 121.29 0 123.15 342.72 ;
      RECT 118.77 0 120.63 342.72 ;
      RECT 113.73 0 118.11 342.72 ;
      RECT 111.21 0 113.07 342.72 ;
      RECT 108.69 0 110.55 342.72 ;
      RECT 98.61 0 108.03 342.72 ;
      RECT 86.01 0 95.43 342.72 ;
      RECT 73.41 0 82.83 342.72 ;
      RECT 60.81 0 70.23 342.72 ;
      RECT 48.21 0 57.63 342.72 ;
      RECT 35.61 0 45.03 342.72 ;
      RECT 23.01 0 32.43 342.72 ;
      RECT 10.41 0 19.83 342.72 ;
      RECT 0 0 7.23 342.72 ;
    LAYER m1 SPACING 0.18 ;
      RECT 0 0 302.4 342.72 ;
  END
END s10hv_1prf_w1024x16b1c08_ulm

END LIBRARY

